`ifndef ALU_REGS_PKG__SV
`define ALU_REGS_PKG__SV

  package alu_regs_pkg;

    // Import UVM
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // Include Reg Model UVCs

  endpackage

`endif

//End of alu_regs_pkg
