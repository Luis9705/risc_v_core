`ifndef CORE_RV32I_REGS_PKG__SV
`define CORE_RV32I_REGS_PKG__SV

  package core_rv32i_regs_pkg;

    // Import UVM
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // Include Reg Model UVCs

  endpackage

`endif

//End of core_rv32i_regs_pkg
