`ifndef COMMON_PKG_SV
`define COMMON_PKG_SV

package common_pkg;

    `define DATA_WIDTH 32
    typedef logic [`DATA_WIDTH-1:0]                data_t;
    
endpackage

`endif

//End of common_pkg