`ifndef REG_FILE_REGS_PKG__SV
`define REG_FILE_REGS_PKG__SV

  package reg_file_regs_pkg;

    // Import UVM
    import uvm_pkg::*;
    `include "uvm_macros.svh"

    // Include Reg Model UVCs

  endpackage

`endif

//End of reg_file_regs_pkg
